`timescale 1 ns / 10 ps

module AvgPoolMulti_tb2 ();
 
reg clk,reset;
reg [16*10*10*16-1:0] inAvg;
wire [16*5*5*16-1:0] outAvg;

localparam PERIOD = 100;

integer i;

always
	#(PERIOD/2) clk = ~clk;
	
initial begin
    #0
    clk = 1'b0;
	  reset = 1;
    inAvg = 25600'h33503a603dd33eb03f0c3e9c3d113b803bb93ac739043c633b90390b3498341ea6a837723b413c8a3a5e36272ad9b554bc5ab8c5a06036bc3b423c9c3628b1b6b4a5b8fdbbb8292839bf38c63a693b0db28bb52f2dd4346838c13d7b3b08361d3661369fb5deb33039f83e3a3f023b8831f731082fcb29c836823c223fc5403e3d8c37ec2e85a7a9b13ca51e383f3c533db33de439512a98b463b4e01e1834edb859b77eb7efb5feb8cebab9b8a52dae366a301dbba9bd1abdc2bcdbbb56b492358935f42e11a4fd39e73eaa416d41b8418c3fd63cbe356f2ffa2c9d3d7f3fe73ec838e52e70b0a8ac67b26d2d0c341c3d9e39fcb5e9beacc082bf3fbc95b8e9b00eab9e39aab7bfbdbec0f0c15ac08bbde0bb62b68bb652b512bd11bf1ac08abf65bc09ba43ba00b8edbafbb81abb93bae4affb3a1f350eb91ebbcabd52bc983ade3d0b3d9c3e0e3c9bad10bd21be4ebd9ebbe73bb83da13acb2e17ba05bde4be55bcfabcb4b9fabc19bc10bcd3bdb1bd93bd35bcc0bc7cba05b545bf81c092c0cec058bf3bbe82bd2dba28b4fdac06ae8db9dbc0a5c440c50ec4b3c266bf54bcc9b8cab9a3c04cc3c7c46dc3b3c24dc024bac0b9b3b877be70c1d3c1f8bfbcbc9abb66b8ddb6d5b95bb919c015c03cbc8eae6430c9b503ba7ebc0bbac8b7d9bd48bbcab6eb342c363ab775be27bec5bbafaddfba19b861b7fd2c8ab7d6bf1dc042bdfeb7a73707bf10bf15bef6c00fc20dc142be58b9642bdd39b6c213c396c403c3f5c222bd8bb61aacda35de3930c062c165c00fbc0dace134cf32b7360c38523465b57a30b13c473d893b07385f392138bc342e2945a2a0b084b528a44c368b3c1139273442315d32a2b473b791b62db2b3b1d0b38cb577af6230d0311fb88ab6d32f7538393450b4f3a654393e3a1134f4b89333a43cdb3d3b3653b39033523da53cdd3390abf83d533f5c3ce635262da83a043f453cd6aae339ef40503f7b3c37396438d13c613eba3a6bb62a3abf3fec3e173aa83a9f39a23b603bbf30e0b52f27843503b78fbbc4b6e19f6634d3323badb2ae12b5d1b596bad2bc9fb9fcac3e2fc22a2daa3728e8a93434d634fc34c3343934983065258d28ca26a838653e55412f41e7414a3e84396a3691376338203d34404a40713f9f389db290ba29b87a302535973f053f553d5f352bbb61bbccbb32b8c8ad23342c3e843d2f368ebc27bcdaa58237389dce25e6b0a03c7f380fb68bbaf82f4e3eff3d90308cb7adb9f23a273535361c3bd43fc540ad3c15b607bbd3bac33bae3ccb3f9d40d1403f3d1833adba86bc20b99f3a4039e039923b0d3ab4322cba31bc8eba83b2daac7bb812ba4aba10bc43be02bdd9bad0b28f27acada2b993bd63bf18bf82bd8eb8baad3f295326ad3b783de63e7e3eeb3e083d3a3c39318eb4f8b17d3d123ce73be4367d303e391a3c09375ab12fb3a53c9838e532f0b4c330ec3c113dda3af22d26b4053b2534b3ab6c34c63c0c3d373d723aa7303bb5e43c0c38b038ed3c4e3bf63ba33b70383cb111b6723e7d3e2b3d2c3d093b8139f43a3c35cfb03db4333ff340133da13c413ad3378230ec28f9a8f5b37a3ea33e37384bb097b63db7d6b0f730d1af9db19e3623347db66fbbb6ba1bafd433b02e6faeadafefb0c6b4d5b140340e37d6368630c5ac04ae84a85234e834392cd62ee6343a37f23c0f3c413df33c12316e2760ac7126ecb0ed2dae3382352e3c7f3c472c1fad9830feb138b204b23e2cb1b1de39c93affb0ceaef2352f3492349bb44fb3f5b22e382a3893b1d835cd3bb63c6e382d2a8eac3834ef360f35c6a9503b633eea3f613b6634eb350937243418315db63734a73b273ca83b4135ea313334723338228eb9b8b91db7eea04a2e80ac242c0932e32f05aeb0b9afb936b8a1b808b4a5aa702bac2c9dad02ae5ab5d5b7ecb929b887b510ad0bac63b061ae35a00d3481383a39923aaf37ca3036b50ab437b5dda9a4381439263b223aad31efb264acb336e932da2c9138f43aa43a2226fcb4812d623bce3bf93a072e8c3a40394e2c85b80535573c9d3e983c4039c0a9053a7334e8b55eaa7c3d553d9b3c5d376f308bafa138112e3c26783aaa3da13b4337b6b190b1b030f0348e34e134bf3a1a3aa1347fb45ab870ad6f37303564375138e83ab4350db496b887b5a2362c3971356737343821364db215b8ddb3e03763397f3580345334c535353412307836ac3a8d39833509287ab919b7043b75414b41283d71324cb880b71fb53ab6163c0a424643b441e73dabad62b9f9b881b6a03b0e4159436341f940a23cbd36d62d8babd1b7a3405641ec413f3cd53b463c693ecc3d5535efba473fd43e8a3965bae1b7013cd240ef3eec330fbb793df63888b966bdab35a14062415e3db624a5bacb3ed13cd5371f38b8402f40af3ec8395eb0f0ba1d3ef83eec3e113e9c3ed83c0936dcac59b712b54c40843faf3cf338ec323badafb4d5b702b403adff4247418c3e44387e32e1addeb36ab196adf8a8a1bc3abd98b96c390f3f4a40a140f93f3f3c80307abcfbb56b3d67418a440a4461448d437940683a61b6113cc740c5435e4499445e448d4403417d3cf23a453f8d4104426c4254416a4253425541533e443ba03e99400b3ebf3b4139133fb14187419240193a803d223b2a34dfb01436c43fd141b4419a3f9e3cbb3dbd3c673c553c033e36407f411f40653dee404d418541b041e540a1404240e040983e513a684185440c44bd446642c0420941453ebe3a522d9040e142d343af43fe4389416d3de2387a2b64a72a3c533ff140703e873c3734972c0029e638dd3a4b3eac3de233eabf2ec1cbc230c0c6bedab791381d3ca2b6a5c0a0c40cc477c3a6c16ec015bc9fb150b6b9c027c1d1c254c214c136c08bbe9fbd00bb41bd2dbed4bd20b901b644bac6bcaebc33bdc7be6fb9e22ebc3c583ead3dbc2cbabc9ebd3cbe96bf09b05c3b653dd73f353a24bc07bfe9becbbdbfbd8cb942b4d0bb4fbe42c05bc13bc068bd8dbc5ebaa6c021c1d9c46ac4aac36ac109be50bc47b9a4b669c2a2c3fec4c7c472c20abf2dbc8bb9f3b657ad64b6eebd67beaebab5385e3e96408e3f543c3f34c3bc75bcb02dda406c4372446e4409414e3e613a05bad335b6411a44794528448b42b8404b3eb33cfe360c3fd0435e444943c640fe3f193e4d3eed3ecf3e0840ef425041153baf37be3d693f594013401a3f1b3f4b3e8331b8ba0a356e3ef340a340703f383c85392f349cb8b6b12e3d8c414441133f853c5d3c703ccb3eec3ff5411b425541ec40613ca0345c3ffb41c3444144b84427428140803cc034159b37410542224360436541d23f4b39da2f28a2f68e0cbde6c0b1c219c295c329c2dac111bfa0bdbbba69bfbac0c3c099bf1bbda5b9dba9ba320bb569b82bc001bf53bc522ede3bd23dc13db43c6c3654af70bef0bce7afb33d263f1d3d5e396a38da3a103553bf06bc0c31663a173677b55cba0ba40f3b7d3b48c044bdeab893bbcbbe1bbe72bc0930533dd93d8ec022bf6fbf2ac132c072be29b8d0396c3ec33d04bc55baacbc00be64bde3b85539413dd53d8e39ee35793d613e1e3b943b513e1b3f6a3e363a2730293adf3fe64201428341da40bf3ea839e02fd3a30fbd4cc14bc369c435c4d8c4f1c49dc388c194bd2bc07bc1eec2a0c2b9c3dec414c429c33bc1eebef2c0cdc192c15dc0b3c12dc20fc346c2a4c1c9bff6c0dac0fcbfdcbe4abfccc174c29cc153c0e7c001c0bfc042bfa4c04cc19ac192c105bfffc01bbedfc0f7c1afc336c410c2d1c119c051be94be2fbcbac1d2c3ecc4d7c4b8c30ac13cbf2ebcb6bbb4b9f7c0dbc26cc39ec388c1e7bfd5bc08b943b910b7c1bcbabed0c06bc086be25ba65b881b845b70ab21db506b93cbb11ba46b8d3b861b821b5fcb10ea2f1bb98bbecaf0f3ddc409040903f953f9c3cf337abbc042b98401843ae43de43bd42ab424440413a3bb4464041441544c544a0444f43b34316412d3ac43cb143a9447b43f142fc41af42b2434141133aa740a443a0428740183d7c3e904234433e40933b4040eb41e840733bed39853f5742dc424b40013bdb408540e13e433ae33d5740ca41c440cf3ed13a334085412f406c403840ca4157410140123c72336b417842b34345438342fe41b1405f3c9b32acabb742414410444443854209401c3afc2d0fac45a42e3bd140d942c141263d19b697be34bd5dbc3db5293ff9411d3d78b76cbd0ebaefbb51b55ab8e9b6553fb73adcbaaec008bfe0b916b5912e5eb807bacc3937b805bde6c0e8bfcfb62031acad45ba6cbe32b55fb8ecbd77beb2b51039e13192b99fbd8fbf46ae6b322e2cdb3aa93ed23788bcafbe55be44bd30397f3b9339be379bb8ffc036c079beffbcf6bb1f3c8d3966bc8dc06dc13fc08ebe6fbd17bb77b7a3ac2cb468bd95bf3cbe30bc86bbebba6db6c4b211bc97bc1abc28bb5fbad9bbaab9b1b618b18caaf3;
    #(PERIOD)
	  reset = 0;
    #(17*PERIOD)
    for (i = 16*5*5-1; i >=0; i = i - 1) begin
		  $displayh(outAvg[i*16+:16]);
	  end
    $stop;
end
AvgPoolMulti 
  #(
  .D(16),
  .H(10),
  .W(10)
  )UUT
  (
    .clk(clk),
    .reset(reset),
    .apInput(inAvg),
    .apOutput(outAvg)
  );
  
endmodule
