`timescale 100 ns / 10 ps

module convLayerMulti_tb();
  
reg reset, clk;
reg [1*32*32*16-1:0] image;
reg [6*1*5*5*16-1:0] filters;
wire [6*28*28*16-1:0] outputConv;

localparam PERIOD = 100;

integer i;
integer file;
always
	#(PERIOD/2) clk = ~clk;
	
initial begin
	$dumpfile("convLayerMulti.vcd");
	$dumpvars(0,convLayerMulti_tb);
end
initial begin
file=$fopen("E:/yanjiusheng/study/研一上/机器学习基础/大作业_曲广龙_杨晓龙/source code/verilog/Conv/result_verilog.txt","w");
end

initial begin 
	#0
	clk = 1'b0;
	reset = 1;
	
	 image = 16384'h3b5f3bc03ba83ba83be03b0f3bf83ba03b7f3bd83aef3b2f3be03be03bb83a9f3bd83c003b983b903bc83ba03bd038c53b1f3bd83bc03ba83b673b7f3be83ba83bb03c003b473bb03b6f3aef3b883b903c003b903b6f3b983bc83b903ac73a363b6f3b473bc83bb03bb03b903bc03a363b773be03bd03bb83c003be03c003b573bb83bb03a663ba03bb03b883b903bb03b903a4e3b2f3bb83bc83bf03b473b773be03b0f3bd83b773b5f3b573ba83b983c003ba03b173ab73bd03b773b3f39ae3bc83b1739753adf3bf83be03bc83bc03bd03a973b3f3bc83b7f3bb03bb83bc03bb83b373bb83b883b7f3b373bc83bc83bd83b5f3b173a873bf03ba83c003aaf3bf03ac738d5393d3adf3a873b5f3be03bf03b903b7f3be03b4f3b3f3be03b1f3a7e3b5f3bb83bd83bc03af73bf83b6f3b7f3bc03c003b3f3bf83b673c003b903bb03aaf387c37983905389d3a7e3bf83b5f3bd03b903be03b773b4f3be83ac73a873bf03bd03b773b273a4e3be83b983bc03bd83bd03b573be83b473b4f3a1e3b883b0f389d37c8386437f839553adf3b983bf03be83bb83b903b7f3b573ac73b983c003bb83af73af73a9f3bb83bd03ba83ba03b473b673c003bf83b7739fe3bd83bc8391d38e538dd3854383c391d3b7f3b6f3bd03b673ba03c003b6f3bc83be83b7f3b883b0f3be03be03bb03bb03b903c003bd03bc03b903b4f3b0f3a463b6f3be03b073b073b7738a537b838d539d63bd03b173bb03c003bc83b673ba03b573be03be03b903bb03bd03bb83bb03bd83b0f3c003b983be03bb03bc03bf03b903bd83ba83b773be83b073a36383c392d3bc83bc83b073b173b903bb03c003c003be83b373aef3b883bf03bc83b983bb03c003c003b5f3a8f3b883bb03ba03ba83b883c003b673aff3ba03b7f37a838ad3b3f3be03b073b883bd03bd83b883ba83bb83b773b5f3bb03bc03ba83bd03b673c003b1f3b673a2e3bc03bd03ba83bf83b473bf83b773af73b983b4f376738543acf3b883b7f3c003b173bb83b273b573bc83be83be03bd83b903b7f3be03ba03b6f3a0e3bd83b2f3bf03bc83bc03c003b6f3bd03b673bd83c003aaf370738043b273b773b983b4f39c63bb03b3f3bc03bd83ba03b7f3bb83bb03b983bc03c003b573a5e3c003be83ba83bb03bb03b6f3bc83bc03a0e3a463a6e3945371738853b983b903ba83b4f3a663bd83a973acf3b6f3ba83b883bb03bc83bc03bd83bd83b983b6f3bd83ba83b7f3be03bd03b473bc03b9838f53834383c383c38543a063b903ba03be03bc83bd83ba03a763a463b673bf03bb03bb03bd03bb83ba03b903b983bf03bb83b573bc03bc03bb83be83b883b7739553874383c3895394d3b4f3b573bb83be83b673be03b1f3b983bb03c003bb83b1f3b773bf03b903ae73bd83b773bd83be83b673c003b273b273c003aff3bb839ce382438a5386c38ad3abf3b983bb039653b573b773b2f3bd03bd03c003a5e38743b4f3b5f3be0394d3b4f3c003b1f3bb03bf83be03b473b2f3ba83bb03bc83ba039753abf38f5380c38cd3b373b983ac73b573bb83ba03b7f3bf83b173a5e3acf3c00399e3aaf3bb83bd03b2f39de3b473be03b903b773c003b773bc83b0f3b4f39e63bd03a76389538343b573b983bb03a873b6f3be83b5f3b4f3bf03b6f3b273bd83af73bc03bd83bf83ba03aef3bb83bd83bc83ba83ba03aff3b903bb03b3f3b5f3bf83bd038bd386c3acf3b7f3ba839f63b0f3bb03b373b6f3bc83b173b473bd83bb83bd83ba03adf3b673bc83be83b983bc03be03b7f3b273bc03c003b773bb83b3f3ba03885389539ee3bd03be03b1f3bd83bd03b903bc03bb83b5f3bf83be83b883ba83c003b883b4f3bc03bc83b773b4f3bb03c003b773bb83b903bc83aff3ae73aa738a5381439053af73a8f3aff3b4f3adf3af73acf3b373b273ad73ab73b1f3b273acf3b3f3af73b2f3a8f3acf3ae73ad73adf3b4f3abf3a363bc03a9f3adf398e384438dd3a973b3f3a763b573b5f3b1f3b573bc03b0f3b373b5f3b983b5f3b2f3aff3aff3b373bb83af73bd83bf03b903bb83bb8397d380c3935389d393d386c37d8383c3b373adf3a3e3b0f3ae73aaf3ab73ac73a9f3b2f3ab73acf3abf3abf3a363b3f3aa73b273aff3ba03a4e39fe3bc83aa73a56375736b7374736c7366637d835a6399639f639553a06398638c539be39d639de39ce39ae39b639de39d639ae39d639fe39b639ce3aaf3b473b5f3b983a363a163854386c3864386439053a5e3aaf3bd03bf03b773bb03bf03be03c003bc03bc83bd03bd83bd83bd03bd03bd03bb83b6f3bc03c003bf83bd83bf03bd03b883ae7398e39f639e63a5e3b1f3c003bc83b903be03be03b7f3be83bd83aa73b473b4f3b883bd83bd83ba83bb03be83c003bf03aa73a6e3b983b373aaf3bd83b983b773b5f3c003b903bd83b983b273bb83b473bb83bf03b7f3bb83b6739f63b4f3b473b883be03bc03b4f3b3f3b983b5f3bc83ac73a663b5f3aff3a7e3bb03be83be83bb83b1f39fe3b2f3c003c003be03bc83bc83bb83bc03bf83bf03b983b903b6f3b903bb83b673abf3a973ad73b883b5f3c003ba0399e3a063bb03bb83b3f3b903be83b883aa73bc83bc03b673b773bb03b883b5f3b7f3b883b903be83bf03be03bf03c003bd03b673b473b673ba83b773bf83b0f393539ee3bc03bc03c003bb03ba83b7f3b273c003bb03ba83bc03bc03be83bf83bd03ba83ba83ba83b883b903b983ba83ba83ba83ba83ba83b6f3bf03be03ba03bd03bd03ba03ba83b883b673bd83bf83b673bc03b3f3c003be83b4f3b983be83b773ba03c003b983bc03bc83bb83ba03ba83bc83bc83ba03bc83b673b983bd83ba83ba83bd03b98;
	 filters[0*5*5*16+:5*5*16] = 400'h2f102cbe28223072b0f4adaf29cb264bab9433cf2dccad87b05f2c8532f1b17a9e72aeadadd428472cf3ade23091b34db1db;
  	 filters[1*5*5*16+:5*5*16] = 400'h282c2cd53092a88bae7621c4310031832a6b32edab0b2ffdac9831c129a3ad1ea991b3a8ad542b2bb28ab3bb2ff9b253af98;
	 filters[2*5*5*16+:5*5*16] = 400'h2f22b0e3ab9ab09d27c431b32601a9c631402cc530f4ac87ac47acd5ad17ae5eb28530ba2fc6ae07317fa47e302a3152adda;
	 filters[3*5*5*16+:5*5*16] = 400'haf1a2d9831bdb088ad462f30acc9aac22c08aeb12fd1afa1af142f7ead63b224b23130f2adf1abde302ca9edae1db0d8b015;
	 filters[4*5*5*16+:5*5*16] = 400'h9cefa80c2ce530a1afbcac1eac24b1b6ac3e31a1a74aaf8031bc2c742992af4da7ceb2b4b212303ba05aaea930c33064b258;
	 filters[5*5*5*16+:5*5*16] = 400'haa3329d2ab9120b631d0afbeb112b14e2f83ae3fb05db1a0321caf87b110b12431b2ae3c2e8aae3aa43a30acb1102f4e226b;
	#(PERIOD)

	reset = 0;

	
	#(7*1457*PERIOD)
	for (i = 6*28*28-1; i >=0; i = i - 1) begin
		$displayh(outputConv[i*16+:16]);
		$fwrite(file,"%h",outputConv[i*16+:16]);
		$fwrite(file,"\n");
	end
	$fclose(file);
	
	$finish;
end

convLayerMulti UUT
(
	.clk(clk),
	.reset(reset),
	.image(image),
	.filters(filters),
	.outputConv(outputConv)
);

endmodule
