`timescale 1 ns / 10 ps

module AvgPoolSingle_TB ();
  
reg [28*28*16-1:0] inAvg;
wire [14*14*16-1:0] outAvg;
initial begin
  $dumpfile("avgpoolsingle.vcd");
  $dumpvars(0,AvgPoolSingle_TB);
end
initial begin
    #0
    inAvg = 12544'h4000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200;
    #10
    $stop;
end
avgPoolSingle UUT
  (
    .aPoolIn(inAvg),
    .aPoolOut(outAvg)
  );
endmodule
    